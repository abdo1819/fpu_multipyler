module number();

endmodule